`timescale 1ns/1ps

module bfp (
    input        clk,
    input        rst_n,
    input [63:0] key_in,        // ---- FIXED 64-bit KEY ----
    input        start_encrypt,
    input [63:0] pt_in,
    output reg [63:0] ct_out,
    output reg   done_encrypt
);
    
    integer i, idx;
    
   (* keep = "true" *) wire [31:0] P [0:17];
    
    
        assign P[0]  = 32'h243F6A88; assign P[1]  = 32'h85A308D3; assign P[2]  = 32'h13198A2E; assign P[3]  = 32'h03707344;
        assign P[4]  = 32'hA4093822; assign P[5]  = 32'h299F31D0; assign P[6]  = 32'h082EFA98; assign P[7]  = 32'hEC4E6C89;
        assign P[8]  = 32'h452821E6; assign P[9]  = 32'h38D01377; assign P[10] = 32'hBE5466CF; assign P[11] = 32'h34E90C6C;
        assign P[12] = 32'hC0AC29B7; assign P[13] = 32'hC97C50DD; assign P[14] = 32'h3F84D5B5; assign P[15] = 32'hB5470917;
        assign P[16] = 32'h9216D5D9; assign P[17] = 32'h8979FB1B;



      

    // -------------------------------------------------------------
    // S-boxes (1024 entries)
    // -------------------------------------------------------------
   (* keep = "true" *)  wire [31:0] S0 [0:255];
   (* keep = "true" *)  wire [31:0] S1 [0:255];
   (* keep = "true" *)  wire [31:0] S2 [0:255];
   (* keep = "true" *) wire [31:0] S3 [0:255];
    
    
    
    // ---------------- S0 ----------------
    assign S0[0] = 32'hD1310BA6;
    assign S0[1] = 32'h98DFB5AC;
    assign S0[2] = 32'h2FFD72DB;
    assign S0[3] = 32'hD01ADFB7;
    assign S0[4] = 32'hB8E1AFED;
    assign S0[5] = 32'h6A267E96;
    assign S0[6] = 32'hBA7C9045;
    assign S0[7] = 32'hF12C7F99;
    assign S0[8] = 32'h24A19947;
    assign S0[9] = 32'hB3916CF7;
    assign S0[10] = 32'h0801F2E2;
    assign S0[11] = 32'h858EFC16;
    assign S0[12] = 32'h636920D8;
    assign S0[13] = 32'h71574E69;
    assign S0[14] = 32'hA458FEA3;
    assign S0[15] = 32'hF4933D7E;
    assign S0[16] = 32'h0D95748F;
    assign S0[17] = 32'h728EB658;
    assign S0[18] = 32'h718BCD58;
    assign S0[19] = 32'h82154AEE;
    assign S0[20] = 32'h7B54A41D;
    assign S0[21] = 32'hC25A59B5;
    assign S0[22] = 32'h9C30D539;
    assign S0[23] = 32'h2AF26013;
    assign S0[24] = 32'hC5D1B023;
    assign S0[25] = 32'h286085F0;
    assign S0[26] = 32'hCA417918;
    assign S0[27] = 32'hB8DB38EF;
    assign S0[28] = 32'h8E79DCB0;
    assign S0[29] = 32'h603A180E;
    assign S0[30] = 32'h6C9E0E8B;
    assign S0[31] = 32'hB01E8A3E;
    assign S0[32] = 32'hD71577C1;
    assign S0[33] = 32'hBD314B27;
    assign S0[34] = 32'h78AF2FDA;
    assign S0[35] = 32'h55605C60;
    assign S0[36] = 32'hE65525F3;
    assign S0[37] = 32'hAA55AB94;
    assign S0[38] = 32'h57489862;
    assign S0[39] = 32'h63E81440;
    assign S0[40] = 32'h55CA396A;
    assign S0[41] = 32'h2AAB10B6;
    assign S0[42] = 32'hB4CC5C34;
    assign S0[43] = 32'h1141E8CE;
    assign S0[44] = 32'hA15486AF;
    assign S0[45] = 32'h7C72E993;
    assign S0[46] = 32'hB3EE1411;
    assign S0[47] = 32'h636FBC2A;
    assign S0[48] = 32'h2BA9C55D;
    assign S0[49] = 32'h741831F6;
    assign S0[50] = 32'hCE5C3E16;
    assign S0[51] = 32'h9B87931E;
    assign S0[52] = 32'hAFD6BA33;
    assign S0[53] = 32'h6C24CF5C;
    assign S0[54] = 32'h7A325381;
    assign S0[55] = 32'h28958677;
    assign S0[56] = 32'h3B8F4898;
    assign S0[57] = 32'h6B4BB9AF;
    assign S0[58] = 32'hC4BFE81B;
    assign S0[59] = 32'h66282193;
    assign S0[60] = 32'h61D809CC;
    assign S0[61] = 32'hFB21A991;
    assign S0[62] = 32'h487CAC60;
    assign S0[63] = 32'h5DEC8032;
    assign S0[64] = 32'hEF845D5D;
    assign S0[65] = 32'hE98575B1;
    assign S0[66] = 32'hDC262302;
    assign S0[67] = 32'hEB651B88;
    assign S0[68] = 32'h23893E81;
    assign S0[69] = 32'hD396ACC5;
    assign S0[70] = 32'h0F6D6FF3;
    assign S0[71] = 32'h83F44239;
    assign S0[72] = 32'h2E0B4482;
    assign S0[73] = 32'hA4842004;
    assign S0[74] = 32'h69C8F04A;
    assign S0[75] = 32'h9E1F9B5E;
    assign S0[76] = 32'h21C66842;
    assign S0[77] = 32'hF6E96C9A;
    assign S0[78] = 32'h670C9C61;
    assign S0[79] = 32'hABD388F0;
    assign S0[80] = 32'h6A51A0D2;
    assign S0[81] = 32'hD8542F68;
    assign S0[82] = 32'h960FA728;
    assign S0[83] = 32'hAB5133A3;
    assign S0[84] = 32'h6EEF0B6C;
    assign S0[85] = 32'h137A3BE4;
    assign S0[86] = 32'hBA3BF050;
    assign S0[87] = 32'h7EFB2A98;
    assign S0[88] = 32'hA1F1651D;
    assign S0[89] = 32'h39AF0176;
    assign S0[90] = 32'h66CA593E;
    assign S0[91] = 32'h82430E88;
    assign S0[92] = 32'h8CEE8619;
    assign S0[93] = 32'h456F9FB4;
    assign S0[94] = 32'h7D84A5C3;
    assign S0[95] = 32'h3B8B5EBE;
    assign S0[96] = 32'hE06F75D8;
    assign S0[97] = 32'h85C12073;
    assign S0[98] = 32'h401A449F;
    assign S0[99] = 32'h56C16AA6;
    assign S0[100] = 32'h4ED3AA62;
    assign S0[101] = 32'h363F7706;
    assign S0[102] = 32'h1BFEDF72;
    assign S0[103] = 32'h429B023D;
    assign S0[104] = 32'h37D0D724;
    assign S0[105] = 32'hD00A1248;
    assign S0[106] = 32'hDB0FEAD3;
    assign S0[107] = 32'h49F1C09B;
    assign S0[108] = 32'h075372C9;
    assign S0[109] = 32'h80991B7B;
    assign S0[110] = 32'h25D479D8;
    assign S0[111] = 32'hF6E8DEF7;
    assign S0[112] = 32'hE3FE501A;
    assign S0[113] = 32'hB6794C3B;
    assign S0[114] = 32'h976CE0BD;
    assign S0[115] = 32'h04C006BA;
    assign S0[116] = 32'hC1A94FB6;
    assign S0[117] = 32'h409F60C4;
    assign S0[118] = 32'h5E5C9EC2;
    assign S0[119] = 32'h196A2463;
    assign S0[120] = 32'h68FB6FAF;
    assign S0[121] = 32'h3E6C53B5;
    assign S0[122] = 32'h1339B2EB;
    assign S0[123] = 32'h3B52EC6F;
    assign S0[124] = 32'h6DFC511F;
    assign S0[125] = 32'h9B30952C;
    assign S0[126] = 32'hCC814544;
    assign S0[127] = 32'hAF5EBD09;
    assign S0[128] = 32'hBEE3D004;
    assign S0[129] = 32'hDE334AFD;
    assign S0[130] = 32'h660F2807;
    assign S0[131] = 32'h192E4BB3;
    assign S0[132] = 32'hC0CBA857;
    assign S0[133] = 32'h45C8740F;
    assign S0[134] = 32'hD20B5F39;
    assign S0[135] = 32'hB9D3FBDB;
    assign S0[136] = 32'h5579C0BD;
    assign S0[137] = 32'h1A60320A;
    assign S0[138] = 32'hD6A100C6;
    assign S0[139] = 32'h402C7279;
    assign S0[140] = 32'h679F25FE;
    assign S0[141] = 32'hFB1FA3CC;
    assign S0[142] = 32'h8EA5E9F8;
    assign S0[143] = 32'hDB3222F8;
    assign S0[144] = 32'h3C7516DF;
    assign S0[145] = 32'hFD616B15;
    assign S0[146] = 32'h2F501EC8;
    assign S0[147] = 32'hAD0552AB;
    assign S0[148] = 32'h323DB5FA;
    assign S0[149] = 32'hFD238760;
    assign S0[150] = 32'h53317B48;
    assign S0[151] = 32'h3E00DF82;
    assign S0[152] = 32'h9E5C57BB;
    assign S0[153] = 32'hCA6F8CA0;
    assign S0[154] = 32'h1A87562E;
    assign S0[155] = 32'hDF1769DB;
    assign S0[156] = 32'hD542A8F6;
    assign S0[157] = 32'h287EFFC3;
    assign S0[158] = 32'hAC6732C6;
    assign S0[159] = 32'h8C4F5573;
    assign S0[160] = 32'h695B27B0;
    assign S0[161] = 32'hBBCA58C8;
    assign S0[162] = 32'hE1FFA35D;
    assign S0[163] = 32'hB8F011A0;
    assign S0[164] = 32'h10FA3D98;
    assign S0[165] = 32'hFD2183B8;
    assign S0[166] = 32'h4AFCB56C;
    assign S0[167] = 32'h2DD1D35B;
    assign S0[168] = 32'h9A53E479;
    assign S0[169] = 32'hB6F84565;
    assign S0[170] = 32'hD28E49BC;
    assign S0[171] = 32'h4BFB9790;
    assign S0[172] = 32'hE1DDF2DA;
    assign S0[173] = 32'hA4CB7E33;
    assign S0[174] = 32'h62FB1341;
    assign S0[175] = 32'hCEE4C6E8;
    assign S0[176] = 32'hEF20CADA;
    assign S0[177] = 32'h36774C01;
    assign S0[178] = 32'hD07E9EFE;
    assign S0[179] = 32'h2BF11FB4;
    assign S0[180] = 32'h95DBDA4D;
    assign S0[181] = 32'hAE909198;
    assign S0[182] = 32'hEAAD8E71;
    assign S0[183] = 32'h6B93D5A0;
    assign S0[184] = 32'hD08ED1D0;
    assign S0[185] = 32'hAFC725E0;
    assign S0[186] = 32'h8E3C5B2F;
    assign S0[187] = 32'h8E7594B7;
    assign S0[188] = 32'h8FF6E2FB;
    assign S0[189] = 32'hF2122B64;
    assign S0[190] = 32'h8888B812;
    assign S0[191] = 32'h900DF01C;
    assign S0[192] = 32'h4FAD5EA0;
    assign S0[193] = 32'h688FC31C;
    assign S0[194] = 32'hD1CFF191;
    assign S0[195] = 32'hB3A8C1AD;
    assign S0[196] = 32'h2F2F2218;
    assign S0[197] = 32'hBE0E1777;
    assign S0[198] = 32'hEA752DFE;
    assign S0[199] = 32'h8B021FA1;
    assign S0[200] = 32'hE5A0CC0F;
    assign S0[201] = 32'hB56F74E8;
    assign S0[202] = 32'h18ACF3D6;
    assign S0[203] = 32'hCE89E299;
    assign S0[204] = 32'hB4A84FE0;
    assign S0[205] = 32'hFD13E0B7;
    assign S0[206] = 32'h7CC43B81;
    assign S0[207] = 32'hD2ADA8D9;
    assign S0[208] = 32'h165FA266;
    assign S0[209] = 32'h80957705;
    assign S0[210] = 32'h93CC7314;
    assign S0[211] = 32'h211A1477;
    assign S0[212] = 32'hE6AD2065;
    assign S0[213] = 32'h77B5FA86;
    assign S0[214] = 32'hC75442F5;
    assign S0[215] = 32'hFB9D35CF;
    assign S0[216] = 32'hEBCDAF0C;
    assign S0[217] = 32'h7B3E89A0;
    assign S0[218] = 32'hD6411BD3;
    assign S0[219] = 32'hAE1E7E49;
    assign S0[220] = 32'h00250E2D;
    assign S0[221] = 32'h2071B35E;
    assign S0[222] = 32'h226800BB;
    assign S0[223] = 32'h57B8E0AF;
    assign S0[224] = 32'h2464369B;
    assign S0[225] = 32'hF009B91E;
    assign S0[226] = 32'h5563911D;
    assign S0[227] = 32'h59DFA6AA;
    assign S0[228] = 32'h78C14389;
    assign S0[229] = 32'hD95A537F;
    assign S0[230] = 32'h207D5BA2;
    assign S0[231] = 32'h02E5B9C5;
    assign S0[232] = 32'h83260376;
    assign S0[233] = 32'h6295CFA9;
    assign S0[234] = 32'h11C81968;
    assign S0[235] = 32'h4E734A41;
    assign S0[236] = 32'hB3472DCA;
    assign S0[237] = 32'h7B14A94A;
    assign S0[238] = 32'h1B510052;
    assign S0[239] = 32'h9A532915;
    assign S0[240] = 32'hD60F573F;
    assign S0[241] = 32'hBC9BC6E4;
    assign S0[242] = 32'h2B60A476;
    assign S0[243] = 32'h81E67400;
    assign S0[244] = 32'h08BA6FB5;
    assign S0[245] = 32'h571BE91F;
    assign S0[246] = 32'hF296EC6B;
    assign S0[247] = 32'h2A0DD915;
    assign S0[248] = 32'hB6636521;
    assign S0[249] = 32'hE7B9F9B6;
    assign S0[250] = 32'hFF34052E;
    assign S0[251] = 32'hC5855664;
    assign S0[252] = 32'h53B02D5D;
    assign S0[253] = 32'hA99F8FA1;
    assign S0[254] = 32'h08BA4799;
    assign S0[255] = 32'h6E85076A;


    
    
    
// ---------------- S1 ----------------
    assign S1[0] = 32'h4B7A70E9;
    assign S1[1] = 32'hB5B32944;
    assign S1[2] = 32'hDB75092E;
    assign S1[3] = 32'hC4192623;
    assign S1[4] = 32'hAD6EA6B0;
    assign S1[5] = 32'h49A7DF7D;
    assign S1[6] = 32'h9CEE60B8;
    assign S1[7] = 32'h8FEDB266;
    assign S1[8] = 32'hECAA8C71;
    assign S1[9] = 32'h699A17FF;
    assign S1[10] = 32'h5664526C;
    assign S1[11] = 32'hC2B19EE1;
    assign S1[12] = 32'h193602A5;
    assign S1[13] = 32'h75094C29;
    assign S1[14] = 32'hA0591340;
    assign S1[15] = 32'hE4183A3E;
    assign S1[16] = 32'h3F54989A;
    assign S1[17] = 32'h5B429D65;
    assign S1[18] = 32'h6B8FE4D6;
    assign S1[19] = 32'h99F73FD6;
    assign S1[20] = 32'hA1D29C07;
    assign S1[21] = 32'hEFE830F5;
    assign S1[22] = 32'h4D2D38E6;
    assign S1[23] = 32'hF0255DC1;
    assign S1[24] = 32'h4CDD2086;
    assign S1[25] = 32'h8470EB26;
    assign S1[26] = 32'h6382E9C6;
    assign S1[27] = 32'h021ECC5E;
    assign S1[28] = 32'h09686B3F;
    assign S1[29] = 32'h3EBAEFC9;
    assign S1[30] = 32'h3C971814;
    assign S1[31] = 32'h6B6A70A1;
    assign S1[32] = 32'h687F3584;
    assign S1[33] = 32'h52A0E286;
    assign S1[34] = 32'hB79C5305;
    assign S1[35] = 32'hAA500737;
    assign S1[36] = 32'h3E07841C;
    assign S1[37] = 32'h7FDEAE5C;
    assign S1[38] = 32'h8E7D44EC;
    assign S1[39] = 32'h5716F2B8;
    assign S1[40] = 32'hB03ADA37;
    assign S1[41] = 32'hF0500C0D;
    assign S1[42] = 32'hF01C1F04;
    assign S1[43] = 32'h0200B3FF;
    assign S1[44] = 32'hAE0CF51A;
    assign S1[45] = 32'h3CB574B2;
    assign S1[46] = 32'h25837A58;
    assign S1[47] = 32'hDC0921BD;
    assign S1[48] = 32'hD19113F9;
    assign S1[49] = 32'h7CA92FF6;
    assign S1[50] = 32'h94324773;
    assign S1[51] = 32'h22F54701;
    assign S1[52] = 32'h3AE5E581;
    assign S1[53] = 32'h37C2DADC;
    assign S1[54] = 32'hC8B57634;
    assign S1[55] = 32'h9AF3DDA7;
    assign S1[56] = 32'hA9446146;
    assign S1[57] = 32'h0FD0030E;
    assign S1[58] = 32'hECC8C73E;
    assign S1[59] = 32'hA4751E41;
    assign S1[60] = 32'hE238CD99;
    assign S1[61] = 32'h3BEA0E2F;
    assign S1[62] = 32'h3280BBA1;
    assign S1[63] = 32'h183EB331;
    assign S1[64] = 32'h4E548B38;
    assign S1[65] = 32'h4F6DB908;
    assign S1[66] = 32'h6F420D03;
    assign S1[67] = 32'hF60A04BF;
    assign S1[68] = 32'h2CB81290;
    assign S1[69] = 32'h24977C79;
    assign S1[70] = 32'h5679B072;
    assign S1[71] = 32'hBCAF89AF;
    assign S1[72] = 32'hDE9A771F;
    assign S1[73] = 32'hD9930810;
    assign S1[74] = 32'hB38BAE12;
    assign S1[75] = 32'hDCCF3F2E;
    assign S1[76] = 32'h5512721F;
    assign S1[77] = 32'h2E6B7124;
    assign S1[78] = 32'h501ADDE6;
    assign S1[79] = 32'h9F84CD87;
    assign S1[80] = 32'h7A584718;
    assign S1[81] = 32'h7408DA17;
    assign S1[82] = 32'hBC9F9ABC;
    assign S1[83] = 32'hE94B7D8C;
    assign S1[84] = 32'hEC7AEC3A;
    assign S1[85] = 32'hDB851DFA;
    assign S1[86] = 32'h63094366;
    assign S1[87] = 32'hC464C3D2;
    assign S1[88] = 32'hEF1C1847;
    assign S1[89] = 32'h3215D908;
    assign S1[90] = 32'hDD433B37;
    assign S1[91] = 32'h24C2BA16;
    assign S1[92] = 32'h12A14D43;
    assign S1[93] = 32'h2A65C451;
    assign S1[94] = 32'h50940002;
    assign S1[95] = 32'h133AE4DD;
    assign S1[96] = 32'h71DFF89E;
    assign S1[97] = 32'h10314E55;
    assign S1[98] = 32'h81AC77D6;
    assign S1[99] = 32'h5F11199B;
    assign S1[100] = 32'h043556F1;
    assign S1[101] = 32'hD7A3C76B;
    assign S1[102] = 32'h3C11183B;
    assign S1[103] = 32'h5924A509;
    assign S1[104] = 32'hF28FE6ED;
    assign S1[105] = 32'h97F1FBFA;
    assign S1[106] = 32'h9EBABF2C;
    assign S1[107] = 32'h1E153C6E;
    assign S1[108] = 32'h86E34570;
    assign S1[109] = 32'hEAE96FB1;
    assign S1[110] = 32'h860E5E0A;
    assign S1[111] = 32'h5A3E2AB3;
    assign S1[112] = 32'h771FE71C;
    assign S1[113] = 32'h4E3D06FA;
    assign S1[114] = 32'h2965DCB9;
    assign S1[115] = 32'h99E71D0F;
    assign S1[116] = 32'h803E89D6;
    assign S1[117] = 32'h5266C825;
    assign S1[118] = 32'h2E4CC978;
    assign S1[119] = 32'h9C10B36A;
    assign S1[120] = 32'hC6150EBA;
    assign S1[121] = 32'h94E2EA78;
    assign S1[122] = 32'hA5FC3C53;
    assign S1[123] = 32'h1E0A2DF4;
    assign S1[124] = 32'hF2F74EA7;
    assign S1[125] = 32'h361D2B3D;
    assign S1[126] = 32'h1939260F;
    assign S1[127] = 32'h19C27960;
    assign S1[128] = 32'h5223A708;
    assign S1[129] = 32'hF71312B6;
    assign S1[130] = 32'hEBADFE6E;
    assign S1[131] = 32'hEAC31F66;
    assign S1[132] = 32'hE3BC4595;
    assign S1[133] = 32'hA67BC883;
    assign S1[134] = 32'hB17F37D1;
    assign S1[135] = 32'h018CFF28;
    assign S1[136] = 32'hC332DDEF;
    assign S1[137] = 32'hBE6C5AA5;
    assign S1[138] = 32'h65582185;
    assign S1[139] = 32'h68AB9802;
    assign S1[140] = 32'hEECEA50F;
    assign S1[141] = 32'hDB2F953B;
    assign S1[142] = 32'h2AEF7DAD;
    assign S1[143] = 32'h5B6E2F84;
    assign S1[144] = 32'h1521B628;
    assign S1[145] = 32'h29076170;
    assign S1[146] = 32'hECDD4775;
    assign S1[147] = 32'h619F1510;
    assign S1[148] = 32'h13CCA830;
    assign S1[149] = 32'hEB61BD96;
    assign S1[150] = 32'h0334FE1E;
    assign S1[151] = 32'hAA0363CF;
    assign S1[152] = 32'hB5735C90;
    assign S1[153] = 32'h4C70A239;
    assign S1[154] = 32'hD59E9E0B;
    assign S1[155] = 32'hCBAADE14;
    assign S1[156] = 32'hEECC86BC;
    assign S1[157] = 32'h60622CA7;
    assign S1[158] = 32'h9CAB5CAB;
    assign S1[159] = 32'hB2F3846E;
    assign S1[160] = 32'h648B1EAF;
    assign S1[161] = 32'h19BDF0CA;
    assign S1[162] = 32'hA02369B9;
    assign S1[163] = 32'h655ABB50;
    assign S1[164] = 32'h40685A32;
    assign S1[165] = 32'h3C2AB4B3;
    assign S1[166] = 32'h319EE9D5;
    assign S1[167] = 32'hC021B8F7;
    assign S1[168] = 32'h9B540B19;
    assign S1[169] = 32'h875FA099;
    assign S1[170] = 32'h95F7997E;
    assign S1[171] = 32'h623D7DA8;
    assign S1[172] = 32'hF837889A;
    assign S1[173] = 32'h97E32D77;
    assign S1[174] = 32'h11ED935F;
    assign S1[175] = 32'h16681281;
    assign S1[176] = 32'h0E358829;
    assign S1[177] = 32'hC7E61FD6;
    assign S1[178] = 32'h96DEDFA1;
    assign S1[179] = 32'h7858BA99;
    assign S1[180] = 32'h57F584A5;
    assign S1[181] = 32'h1B227263;
    assign S1[182] = 32'h9B83C3FF;
    assign S1[183] = 32'h1AC24696;
    assign S1[184] = 32'hCDB30AEB;
    assign S1[185] = 32'h532E3054;
    assign S1[186] = 32'h8FD948E4;
    assign S1[187] = 32'h6DBC3128;
    assign S1[188] = 32'h58EBF2EF;
    assign S1[189] = 32'h34C6FFEA;
    assign S1[190] = 32'hFE28ED61;
    assign S1[191] = 32'hEE7C3C73;
    assign S1[192] = 32'h5D4A14D9;
    assign S1[193] = 32'hE864B7E3;
    assign S1[194] = 32'h42105D14;
    assign S1[195] = 32'h203E13E0;
    assign S1[196] = 32'h45EEE2B6;
    assign S1[197] = 32'hA3AAABEA;
    assign S1[198] = 32'hDB6C4F15;
    assign S1[199] = 32'hFACB4FD0;
    assign S1[200] = 32'hC742F442;
    assign S1[201] = 32'hEF6ABBB5;
    assign S1[202] = 32'h654F3B1D;
    assign S1[203] = 32'h41CD2105;
    assign S1[204] = 32'hD81E799E;
    assign S1[205] = 32'h86854DC7;
    assign S1[206] = 32'hE44B476A;
    assign S1[207] = 32'h3D816250;
    assign S1[208] = 32'hCF62A1F2;
    assign S1[209] = 32'h5B8D2646;
    assign S1[210] = 32'hFC8883A0;
    assign S1[211] = 32'hC1C7B6A3;
    assign S1[212] = 32'h7F1524C3;
    assign S1[213] = 32'h69CB7492;
    assign S1[214] = 32'h47848A0B;
    assign S1[215] = 32'h5692B285;
    assign S1[216] = 32'h095BBF00;
    assign S1[217] = 32'hAD19489D;
    assign S1[218] = 32'h1462B174;
    assign S1[219] = 32'h23820E00;
    assign S1[220] = 32'h58428D2A;
    assign S1[221] = 32'h0C55F5EA;
    assign S1[222] = 32'h1DADF43E;
    assign S1[223] = 32'h233F7061;
    assign S1[224] = 32'h3372F092;
    assign S1[225] = 32'h8D937E41;
    assign S1[226] = 32'hD65FECF1;
    assign S1[227] = 32'h6C223BDB;
    assign S1[228] = 32'h7CDE3759;
    assign S1[229] = 32'hCBEE7460;
    assign S1[230] = 32'h4085F2A7;
    assign S1[231] = 32'hCE77326E;
    assign S1[232] = 32'hA6078084;
    assign S1[233] = 32'h19F8509E;
    assign S1[234] = 32'hE8EFD855;
    assign S1[235] = 32'h61D99735;
    assign S1[236] = 32'hA969A7AA;
    assign S1[237] = 32'hC50C06C2;
    assign S1[238] = 32'h5A04ABFC;
    assign S1[239] = 32'h800BCADC;
    assign S1[240] = 32'h9E447A2E;
    assign S1[241] = 32'hC3453484;
    assign S1[242] = 32'hFDD56705;
    assign S1[243] = 32'h0E1E9EC9;
    assign S1[244] = 32'hDB73DBD3;
    assign S1[245] = 32'h105588CD;
    assign S1[246] = 32'h675FDA79;
    assign S1[247] = 32'hE3674340;
    assign S1[248] = 32'hC5C43465;
    assign S1[249] = 32'h713E38D8;
    assign S1[250] = 32'h3D28F89E;
    assign S1[251] = 32'hF16DFF20;
    assign S1[252] = 32'h153E21E7;
    assign S1[253] = 32'h8FB03D4A;
    assign S1[254] = 32'hE6E39F2B;
    assign S1[255] = 32'hDB83ADF7;





// ---------------- S2 ----------------
 
    assign S2[0] = 32'hE93D5A68;
    assign S2[1] = 32'h948140F7;
    assign S2[2] = 32'hF64C261C;
    assign S2[3] = 32'h94692934;
    assign S2[4] = 32'h411520F7;
    assign S2[5] = 32'h7602D4F7;
    assign S2[6] = 32'hBCF46B2E;
    assign S2[7] = 32'hD4A20068;
    assign S2[8] = 32'hD4082471;
    assign S2[9] = 32'h3320F46A;
    assign S2[10] = 32'h43B7D4B7;
    assign S2[11] = 32'h500061AF;
    assign S2[12] = 32'h1E39F62E;
    assign S2[13] = 32'h97244546;
    assign S2[14] = 32'h14214F74;
    assign S2[15] = 32'hBF8B8840;
    assign S2[16] = 32'h4D95FC1D;
    assign S2[17] = 32'h96B591AF;
    assign S2[18] = 32'h70F4DDD3;
    assign S2[19] = 32'h66A02F45;
    assign S2[20] = 32'hBFBC09EC;
    assign S2[21] = 32'h03BD9785;
    assign S2[22] = 32'h7FAC6DD0;
    assign S2[23] = 32'h31CB8504;
    assign S2[24] = 32'h96EB27B3;
    assign S2[25] = 32'h55FD3941;
    assign S2[26] = 32'hDA2547E6;
    assign S2[27] = 32'hABCA0A9A;
    assign S2[28] = 32'h28507825;
    assign S2[29] = 32'h530429F4;
    assign S2[30] = 32'h0A2C86DA;
    assign S2[31] = 32'hE9B66DFB;
    assign S2[32] = 32'h68DC1462;
    assign S2[33] = 32'hD7486900;
    assign S2[34] = 32'h680EC0A4;
    assign S2[35] = 32'h27A18DEE;
    assign S2[36] = 32'h4F3FFEA2;
    assign S2[37] = 32'hE887AD8C;
    assign S2[38] = 32'hB58CE006;
    assign S2[39] = 32'h7AF4D6B6;
    assign S2[40] = 32'hAACE1E7C;
    assign S2[41] = 32'hD3375FEC;
    assign S2[42] = 32'hCE78A399;
    assign S2[43] = 32'h406B2A42;
    assign S2[44] = 32'h20FE9E35;
    assign S2[45] = 32'hD9F385B9;
    assign S2[46] = 32'hEE39D7AB;
    assign S2[47] = 32'h3B124E8B;
    assign S2[48] = 32'h1DC9FAF7;
    assign S2[49] = 32'h4B6D1856;
    assign S2[50] = 32'h26A36631;
    assign S2[51] = 32'hEAE397B2;
    assign S2[52] = 32'h3A6EFA74;
    assign S2[53] = 32'hDD5B4332;
    assign S2[54] = 32'h6841E7F7;
    assign S2[55] = 32'hCA7820FB;
    assign S2[56] = 32'hFB0AF54E;
    assign S2[57] = 32'hD8FEB397;
    assign S2[58] = 32'h454056AC;
    assign S2[59] = 32'hBA489527;
    assign S2[60] = 32'h55533A3A;
    assign S2[61] = 32'h20838D87;
    assign S2[62] = 32'hFE6BA9B7;
    assign S2[63] = 32'hD096954B;
    assign S2[64] = 32'h55A867BC;
    assign S2[65] = 32'hA1159A58;
    assign S2[66] = 32'hCCA92963;
    assign S2[67] = 32'h99E1DB33;
    assign S2[68] = 32'hA62A4A56;
    assign S2[69] = 32'h3F3125F9;
    assign S2[70] = 32'h5EF47E1C;
    assign S2[71] = 32'h9029317C;
    assign S2[72] = 32'hFDF8E802;
    assign S2[73] = 32'h04272F70;
    assign S2[74] = 32'h80BB155C;
    assign S2[75] = 32'h05282CE3;
    assign S2[76] = 32'h95C11548;
    assign S2[77] = 32'hE4C66D22;
    assign S2[78] = 32'h48C1133F;
    assign S2[79] = 32'hC70F86DC;
    assign S2[80] = 32'h07F9C9EE;
    assign S2[81] = 32'h41041F0F;
    assign S2[82] = 32'h404779A4;
    assign S2[83] = 32'h5D886E17;
    assign S2[84] = 32'h325F51EB;
    assign S2[85] = 32'hD59BC0D1;
    assign S2[86] = 32'hF2BCC18F;
    assign S2[87] = 32'h41113564;
    assign S2[88] = 32'h257B7834;
    assign S2[89] = 32'h602A9C60;
    assign S2[90] = 32'hDFF8E8A3;
    assign S2[91] = 32'h1F636C1B;
    assign S2[92] = 32'h0E12B4C2;
    assign S2[93] = 32'h02E1329E;
    assign S2[94] = 32'hAF664FD1;
    assign S2[95] = 32'hCAD18115;
    assign S2[96] = 32'h6B2395E0;
    assign S2[97] = 32'h333E92E1;
    assign S2[98] = 32'h3B240B62;
    assign S2[99] = 32'hEEBEB922;
    assign S2[100] = 32'h85B2A20E;
    assign S2[101] = 32'hE6BA0D99;
    assign S2[102] = 32'hDE720C8C;
    assign S2[103] = 32'h2DA2F728;
    assign S2[104] = 32'hD0127845;
    assign S2[105] = 32'h95B794FD;
    assign S2[106] = 32'h647D0862;
    assign S2[107] = 32'hE7CCF5F0;
    assign S2[108] = 32'h5449A36F;
    assign S2[109] = 32'h877D48FA;
    assign S2[110] = 32'hC39DFD27;
    assign S2[111] = 32'hF33E8D1E;
    assign S2[112] = 32'h0A476341;
    assign S2[113] = 32'h992EFF74;
    assign S2[114] = 32'h3A6F6EAB;
    assign S2[115] = 32'hF4F8FD37;
    assign S2[116] = 32'hA812DC60;
    assign S2[117] = 32'hA1EBDDF8;
    assign S2[118] = 32'h991BE14C;
    assign S2[119] = 32'hDB6E6B0D;
    assign S2[120] = 32'hC67B5510;
    assign S2[121] = 32'h6D672C37;
    assign S2[122] = 32'h2765D43B;
    assign S2[123] = 32'hDCD0E804;
    assign S2[124] = 32'hF1290DC7;
    assign S2[125] = 32'hCC00FFA3;
    assign S2[126] = 32'hB5390F92;
    assign S2[127] = 32'h690FED0B;
    assign S2[128] = 32'h667B9FFB;
    assign S2[129] = 32'hCEDB7D9C;
    assign S2[130] = 32'hA091CF0B;
    assign S2[131] = 32'hD9155EA3;
    assign S2[132] = 32'hBB132F88;
    assign S2[133] = 32'h515BAD24;
    assign S2[134] = 32'h7B9479BF;
    assign S2[135] = 32'h763BD6EB;
    assign S2[136] = 32'h37392EB3;
    assign S2[137] = 32'hCC115979;
    assign S2[138] = 32'h8026E297;
    assign S2[139] = 32'hF42E312D;
    assign S2[140] = 32'h6842ADA7;
    assign S2[141] = 32'hC66A2B3B;
    assign S2[142] = 32'h12754CCC;
    assign S2[143] = 32'h782EF11C;
    assign S2[144] = 32'h6A124237;
    assign S2[145] = 32'hB79251E7;
    assign S2[146] = 32'h06A1BBE6;
    assign S2[147] = 32'h4BFB6350;
    assign S2[148] = 32'h1A6B1018;
    assign S2[149] = 32'h11CAEDFA;
    assign S2[150] = 32'h3D25BDD8;
    assign S2[151] = 32'hE2E1C3C9;
    assign S2[152] = 32'h44421659;
    assign S2[153] = 32'h0A121386;
    assign S2[154] = 32'hD90CEC6E;
    assign S2[155] = 32'hD5ABEA2A;
    assign S2[156] = 32'h64AF674E;
    assign S2[157] = 32'hDA86A85F;
    assign S2[158] = 32'hBEBFE988;
    assign S2[159] = 32'h64E4C3FE;
    assign S2[160] = 32'h9DBC8057;
    assign S2[161] = 32'hF0F7C086;
    assign S2[162] = 32'h60787BF8;
    assign S2[163] = 32'h6003604D;
    assign S2[164] = 32'hD1FD8346;
    assign S2[165] = 32'hF6381FB0;
    assign S2[166] = 32'h7745AE04;
    assign S2[167] = 32'hD736FCCC;
    assign S2[168] = 32'h83426B33;
    assign S2[169] = 32'hF01EAB71;
    assign S2[170] = 32'hB0804187;
    assign S2[171] = 32'h3C005E5F;
    assign S2[172] = 32'h77A057BE;
    assign S2[173] = 32'hBDE8AE24;
    assign S2[174] = 32'h55464299;
    assign S2[175] = 32'hBF582E61;
    assign S2[176] = 32'h4E58F48F;
    assign S2[177] = 32'hF2DDFDA2;
    assign S2[178] = 32'hF474EF38;
    assign S2[179] = 32'h8789BDC2;
    assign S2[180] = 32'h5366F9C3;
    assign S2[181] = 32'hC8B38E74;
    assign S2[182] = 32'hB475F255;
    assign S2[183] = 32'h46FCD9B9;
    assign S2[184] = 32'h7AEB2661;
    assign S2[185] = 32'h8B1DDF84;
    assign S2[186] = 32'h846A0E79;
    assign S2[187] = 32'h915F95E2;
    assign S2[188] = 32'h466E598E;
    assign S2[189] = 32'h20B45770;
    assign S2[190] = 32'h8CD55591;
    assign S2[191] = 32'hC902DE4C;
    assign S2[192] = 32'hB90BACE1;
    assign S2[193] = 32'hBB8205D0;
    assign S2[194] = 32'h11A86248;
    assign S2[195] = 32'h7574A99E;
    assign S2[196] = 32'hB77F19B6;
    assign S2[197] = 32'hE0A9DC09;
    assign S2[198] = 32'h662D09A1;
    assign S2[199] = 32'hC4324633;
    assign S2[200] = 32'hE85A1F02;
    assign S2[201] = 32'h09F0BE8C;
    assign S2[202] = 32'h4A99A025;
    assign S2[203] = 32'h1D6EFE10;
    assign S2[204] = 32'h1AB93D1D;
    assign S2[205] = 32'h0BA5A4DF;
    assign S2[206] = 32'hA186F20F;
    assign S2[207] = 32'h2868F169;
    assign S2[208] = 32'hDCB7DA83;
    assign S2[209] = 32'h573906FE;
    assign S2[210] = 32'hA1E2CE9B;
    assign S2[211] = 32'h4FCD7F52;
    assign S2[212] = 32'h50115E01;
    assign S2[213] = 32'hA70683FA;
    assign S2[214] = 32'hA002B5C4;
    assign S2[215] = 32'h0DE6D027;
    assign S2[216] = 32'h9AF88C27;
    assign S2[217] = 32'h773F8641;
    assign S2[218] = 32'hC3604C06;
    assign S2[219] = 32'h61A806B5;
    assign S2[220] = 32'hF0177A28;
    assign S2[221] = 32'hC0F586E0;
    assign S2[222] = 32'h006058AA;
    assign S2[223] = 32'h30DC7D62;
    assign S2[224] = 32'h11E69ED7;
    assign S2[225] = 32'h2338EA63;
    assign S2[226] = 32'h53C2DD94;
    assign S2[227] = 32'hC2C21634;
    assign S2[228] = 32'hBBCBEE56;
    assign S2[229] = 32'h90BCB6DE;
    assign S2[230] = 32'hEBFC7DA1;
    assign S2[231] = 32'hCE591D76;
    assign S2[232] = 32'h6F05E409;
    assign S2[233] = 32'h4B7C0188;
    assign S2[234] = 32'h39720A3D;
    assign S2[235] = 32'h7C927C24;
    assign S2[236] = 32'h86E3725F;
    assign S2[237] = 32'h724D9DB9;
    assign S2[238] = 32'h1AC15BB4;
    assign S2[239] = 32'hD39EB8FC;
    assign S2[240] = 32'hED545578;
    assign S2[241] = 32'h08FCA5B5;
    assign S2[242] = 32'hD83D7CD3;
    assign S2[243] = 32'h4DAD0FC4;
    assign S2[244] = 32'h1E50EF5E;
    assign S2[245] = 32'hB161E6F8;
    assign S2[246] = 32'hA28514D9;
    assign S2[247] = 32'h6C51133C;
    assign S2[248] = 32'h6FD5C7E7;
    assign S2[249] = 32'h56E14EC4;
    assign S2[250] = 32'h362ABFCE;
    assign S2[251] = 32'hDDC6C837;
    assign S2[252] = 32'hD79A3234;
    assign S2[253] = 32'h92638212;
    assign S2[254] = 32'h670EFA8E;
    assign S2[255] = 32'h406000E0;



// ---------------- S3 ----------------
    assign S3[0] = 32'h3A39CE37;
    assign S3[1] = 32'hD3FAF5CF;
    assign S3[2] = 32'hABC27737;
    assign S3[3] = 32'h5AC52D1B;
    assign S3[4] = 32'h5CB0679E;
    assign S3[5] = 32'h4FA33742;
    assign S3[6] = 32'hD3822740;
    assign S3[7] = 32'h99BC9BBE;
    assign S3[8] = 32'hD5118E9D;
    assign S3[9] = 32'hBF0F7315;
    assign S3[10] = 32'hD62D1C7E;
    assign S3[11] = 32'hC700C47B;
    assign S3[12] = 32'hB78C1B6B;
    assign S3[13] = 32'h21A19045;
    assign S3[14] = 32'hB26EB1BE;
    assign S3[15] = 32'h6A366EB4;
    assign S3[16] = 32'h5748AB2F;
    assign S3[17] = 32'hBC946E79;
    assign S3[18] = 32'hC6A376D2;
    assign S3[19] = 32'h6549C2C8;
    assign S3[20] = 32'h530FF8EE;
    assign S3[21] = 32'h468DDE7D;
    assign S3[22] = 32'hD5730A1D;
    assign S3[23] = 32'h4CD04DC6;
    assign S3[24] = 32'h2939BBDB;
    assign S3[25] = 32'hA9BA4650;
    assign S3[26] = 32'hAC9526E8;
    assign S3[27] = 32'hBE5EE304;
    assign S3[28] = 32'hA1FAD5F0;
    assign S3[29] = 32'h6A2D519A;
    assign S3[30] = 32'h63EF8CE2;
    assign S3[31] = 32'h9A86EE22;
    assign S3[32] = 32'hC089C2B8;
    assign S3[33] = 32'h43242EF6;
    assign S3[34] = 32'hA51E03AA;
    assign S3[35] = 32'h9CF2D0A4;
    assign S3[36] = 32'h83C061BA;
    assign S3[37] = 32'h9BE96A4D;
    assign S3[38] = 32'h8FE51550;
    assign S3[39] = 32'hBA645BD6;
    assign S3[40] = 32'h2826A2F9;
    assign S3[41] = 32'hA73A3AE1;
    assign S3[42] = 32'h4BA99586;
    assign S3[43] = 32'hEF5562E9;
    assign S3[44] = 32'hC72FEFD3;
    assign S3[45] = 32'hF752F7DA;
    assign S3[46] = 32'h3F046F69;
    assign S3[47] = 32'h77FA0A59;
    assign S3[48] = 32'h80E4A915;
    assign S3[49] = 32'h87B08601;
    assign S3[50] = 32'h9B09E6AD;
    assign S3[51] = 32'h3B3EE593;
    assign S3[52] = 32'hE990FD5A;
    assign S3[53] = 32'h9E34D797;
    assign S3[54] = 32'h2CF0B7D9;
    assign S3[55] = 32'h022B8B51;
    assign S3[56] = 32'h96D5AC3A;
    assign S3[57] = 32'h017DA67D;
    assign S3[58] = 32'hD1CF3ED6;
    assign S3[59] = 32'h7C7D2D28;
    assign S3[60] = 32'h1F9F25CF;
    assign S3[61] = 32'hADF2B89B;
    assign S3[62] = 32'h5AD6B472;
    assign S3[63] = 32'h5A88F54C;
    assign S3[64] = 32'hE029AC71;
    assign S3[65] = 32'hE019A5E6;
    assign S3[66] = 32'h47B0ACFD;
    assign S3[67] = 32'hED93FA9B;
    assign S3[68] = 32'hE8D3C48D;
    assign S3[69] = 32'h283B57CC;
    assign S3[70] = 32'hF8D56629;
    assign S3[71] = 32'h79132E28;
    assign S3[72] = 32'h785F0191;
    assign S3[73] = 32'hED756055;
    assign S3[74] = 32'hF7960E44;
    assign S3[75] = 32'hE3D35E8C;
    assign S3[76] = 32'h15056DD4;
    assign S3[77] = 32'h88F46DBA;
    assign S3[78] = 32'h03A16125;
    assign S3[79] = 32'h0564F0BD;
    assign S3[80] = 32'hC3EB9E15;
    assign S3[81] = 32'h3C9057A2;
    assign S3[82] = 32'h97271AEC;
    assign S3[83] = 32'hA93A072A;
    assign S3[84] = 32'h1B3F6D9B;
    assign S3[85] = 32'h1E6321F5;
    assign S3[86] = 32'hF59C66FB;
    assign S3[87] = 32'h26DCF319;
    assign S3[88] = 32'h7533D928;
    assign S3[89] = 32'hB155FDF5;
    assign S3[90] = 32'h03563482;
    assign S3[91] = 32'h8ABA3CBB;
    assign S3[92] = 32'h28517711;
    assign S3[93] = 32'hC20AD9F8;
    assign S3[94] = 32'hABCC5167;
    assign S3[95] = 32'hCCAD925F;
    assign S3[96] = 32'h4DE81751;
    assign S3[97] = 32'h3830DC8E;
    assign S3[98] = 32'h379D5862;
    assign S3[99] = 32'h9320F991;
    assign S3[100] = 32'hEA7A90C2;
    assign S3[101] = 32'hFB3E7BCE;
    assign S3[102] = 32'h5121CE64;
    assign S3[103] = 32'h774FBE32;
    assign S3[104] = 32'hA8B6E37E;
    assign S3[105] = 32'hC3293D46;
    assign S3[106] = 32'h48DE5369;
    assign S3[107] = 32'h6413E680;
    assign S3[108] = 32'hA2AE0810;
    assign S3[109] = 32'hDD6DB224;
    assign S3[110] = 32'h69852DFD;
    assign S3[111] = 32'h09072166;
    assign S3[112] = 32'hB39A460A;
    assign S3[113] = 32'h6445C0DD;
    assign S3[114] = 32'h586CDECF;
    assign S3[115] = 32'h1C20C8AE;
    assign S3[116] = 32'h5BBEF7DD;
    assign S3[117] = 32'h1B588D40;
    assign S3[118] = 32'hCCD2017F;
    assign S3[119] = 32'h6BB4E3BB;
    assign S3[120] = 32'hDDA26A7E;
    assign S3[121] = 32'h3A59FF45;
    assign S3[122] = 32'h3E350A44;
    assign S3[123] = 32'hBCB4CDD5;
    assign S3[124] = 32'h72Eacea8;
    assign S3[125] = 32'hFA6484BB;
    assign S3[126] = 32'h8D6612AE;
    assign S3[127] = 32'hBF3C6F47;
    assign S3[128] = 32'hD29BE463;
    assign S3[129] = 32'h542F5D9E;
    assign S3[130] = 32'hAEC2771B;
    assign S3[131] = 32'hF64E6370;
    assign S3[132] = 32'h740E0D8D;
    assign S3[133] = 32'hE75B1357;
    assign S3[134] = 32'hF8721671;
    assign S3[135] = 32'hAF537D5D;
    assign S3[136] = 32'h4040CB08;
    assign S3[137] = 32'h4EB4E2CC;
    assign S3[138] = 32'h34D2466A;
    assign S3[139] = 32'h0115AF84;
    assign S3[140] = 32'hE1B00428;
    assign S3[141] = 32'h95983A1D;
    assign S3[142] = 32'h06B89FB4;
    assign S3[143] = 32'hCE6EA048;
    assign S3[144] = 32'h6F3F3B82;
    assign S3[145] = 32'h3520AB82;
    assign S3[146] = 32'h011A1D4B;
    assign S3[147] = 32'h277227F8;
    assign S3[148] = 32'h611560B1;
    assign S3[149] = 32'hE7933FDC;
    assign S3[150] = 32'hBB3A792B;
    assign S3[151] = 32'h344525BD;
    assign S3[152] = 32'hA08839E1;
    assign S3[153] = 32'h51CE794B;
    assign S3[154] = 32'h2F32C9B7;
    assign S3[155] = 32'hA01FBAC9;
    assign S3[156] = 32'hE01CC87E;
    assign S3[157] = 32'hBCC7D1F6;
    assign S3[158] = 32'hCF0111C3;
    assign S3[159] = 32'hA1E8AAC7;
    assign S3[160] = 32'h1A908749;
    assign S3[161] = 32'hD44FBD9A;
    assign S3[162] = 32'hD0DADECB;
    assign S3[163] = 32'hD50ADA38;
    assign S3[164] = 32'h0339C32A;
    assign S3[165] = 32'hC6913667;
    assign S3[166] = 32'h8DF9317C;
    assign S3[167] = 32'hE0B12B4F;
    assign S3[168] = 32'hF79E59B7;
    assign S3[169] = 32'h43F5BB3A;
    assign S3[170] = 32'hF2D519FF;
    assign S3[171] = 32'h27D9459C;
    assign S3[172] = 32'hBF97222C;
    assign S3[173] = 32'h15E6FC2A;
    assign S3[174] = 32'h0F91FC71;
    assign S3[175] = 32'h9B941525;
    assign S3[176] = 32'hFAE59361;
    assign S3[177] = 32'hCEB69CEB;
    assign S3[178] = 32'hC2A86459;
    assign S3[179] = 32'h12BAA8D1;
    assign S3[180] = 32'hB6C1075E;
    assign S3[181] = 32'hE3056A0C;
    assign S3[182] = 32'h10D25065;
    assign S3[183] = 32'hCB03A442;
    assign S3[184] = 32'hE0EC6E0E;
    assign S3[185] = 32'h1698DB3B;
    assign S3[186] = 32'h4C98A0BE;
    assign S3[187] = 32'h3278E964;
    assign S3[188] = 32'h9F1F9532;
    assign S3[189] = 32'hE0D392DF;
    assign S3[190] = 32'hD3A0342B;
    assign S3[191] = 32'h8971F21E;
    assign S3[192] = 32'h1B0A7441;
    assign S3[193] = 32'h4BA3348C;
    assign S3[194] = 32'hC5BE7120;
    assign S3[195] = 32'hC37632D8;
    assign S3[196] = 32'hDF359F8D;
    assign S3[197] = 32'h9B992F2E;
    assign S3[198] = 32'hE60B6F47;
    assign S3[199] = 32'h0FE3F11D;
    assign S3[200] = 32'hE54CDA54;
    assign S3[201] = 32'h1EDAD891;
    assign S3[202] = 32'hCE6279CF;
    assign S3[203] = 32'hCD3E7E6F;
    assign S3[204] = 32'h1618B166;
    assign S3[205] = 32'hFD2C1D05;
    assign S3[206] = 32'h848FD2C5;
    assign S3[207] = 32'hF6FB2299;
    assign S3[208] = 32'hF523F357;
    assign S3[209] = 32'hA6327623;
    assign S3[210] = 32'h93A83531;
    assign S3[211] = 32'h56CCCD02;
    assign S3[212] = 32'hACF08162;
    assign S3[213] = 32'h5A75EBB5;
    assign S3[214] = 32'h6E163697;
    assign S3[215] = 32'h88D273CC;
    assign S3[216] = 32'hDE966292;
    assign S3[217] = 32'h81B949D0;
    assign S3[218] = 32'h4C50901B;
    assign S3[219] = 32'h71C65614;
    assign S3[220] = 32'hE6C6C7BD;
    assign S3[221] = 32'h327A140A;
    assign S3[222] = 32'h45E1D006;
    assign S3[223] = 32'hC3F27B9A;
    assign S3[224] = 32'hC9AA53FD;
    assign S3[225] = 32'h62A80F00;
    assign S3[226] = 32'hBB25BFE2;
    assign S3[227] = 32'h35BDD2F6;
    assign S3[228] = 32'h71126905;
    assign S3[229] = 32'hB2040222;
    assign S3[230] = 32'hB6CBCF7C;
    assign S3[231] = 32'hCD769C2B;
    assign S3[232] = 32'h53113EC0;
    assign S3[233] = 32'h1640E3D3;
    assign S3[234] = 32'h38ABBD60;
    assign S3[235] = 32'h2547ADF0;
    assign S3[236] = 32'hBA38209C;
    assign S3[237] = 32'hF746CE76;
    assign S3[238] = 32'h77AFA1C5;
    assign S3[239] = 32'h20756060;
    assign S3[240] = 32'h85CBFE4E;
    assign S3[241] = 32'h8AE88DD8;
    assign S3[242] = 32'h7AAAF9B0;
    assign S3[243] = 32'h4CF9AA7E;
    assign S3[244] = 32'h1948C25C;
    assign S3[245] = 32'h02FB8A8C;
    assign S3[246] = 32'h01C36AE4;
    assign S3[247] = 32'hD6EBE1F9;
    assign S3[248] = 32'h90D4F869;
    assign S3[249] = 32'hA65CDEA0;
    assign S3[250] = 32'h3F09252D;
    assign S3[251] = 32'hC208E69F;
    assign S3[252] = 32'hB74E6132;
    assign S3[253] = 32'hCE77E25B;
    assign S3[254] = 32'h578FDFE3;
    assign S3[255] = 32'h3AC372E6;
  function [31:0] F_func;
        input [31:0] x;
        reg [7:0] a,b,c,d;
        reg [31:0] y;
    begin
        a = x[31:24];
        b = x[23:16];
        c = x[15:8];
        d = x[7:0];
        y = S0[a] + S1[b];
        y = y ^  S2[c];
        y = y +  S3[d];
        F_func = y;
    end
    endfunction

    // -------------------------------------------------------------
    // Blowfish Encryption Engine ONLY (16 rounds)
    // -------------------------------------------------------------
    reg        enc_busy;
    reg [4:0]  round;
    reg [31:0] L, R, Ltmp, Rtmp;

    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            enc_busy      <= 0;
            round         <= 0;
            done_encrypt  <= 0;
            ct_out        <= 0;
        end else begin

            // Start only when idle
            if(start_encrypt && !enc_busy) begin
                enc_busy <= 1;
                round    <= 0;
                L <= pt_in[63:32];
                R <= pt_in[31:0];
            end

            // Run 16 rounds
            else if(enc_busy) begin
                if(round < 16) begin
                    Ltmp = L ^  P[round];
                    Rtmp = R ^ F_func(Ltmp);

                    L    <= Rtmp;
                    R    <= Ltmp;
                    round <= round + 1;
                end
                else begin
                    // Final XORs
                    R <= R ^  P[16];
                    L <= L ^  P[17];

                    ct_out <= {L, R};
                    done_encrypt <= 1;
                    enc_busy <= 0;
                end
            end
        end
    end

   
endmodule
